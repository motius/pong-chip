VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pong
  CLASS BLOCK ;
  FOREIGN pong ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN blue[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END blue[0]
  PIN blue[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 374.720 900.000 375.320 ;
    END
  END blue[1]
  PIN blue[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 0.000 675.190 4.000 ;
    END
  END blue[2]
  PIN blue[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.870 0.000 825.150 4.000 ;
    END
  END blue[3]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.870 596.000 825.150 600.000 ;
    END
  END clk
  PIN game_reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END game_reset
  PIN green[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END green[0]
  PIN green[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END green[1]
  PIN green[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.280 4.000 471.880 ;
    END
  END green[2]
  PIN green[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 524.320 900.000 524.920 ;
    END
  END green[3]
  PIN hsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END hsync
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 596.000 25.210 600.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 596.000 525.230 600.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.630 596.000 574.910 600.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 596.000 625.050 600.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 596.000 675.190 600.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 596.000 725.330 600.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.730 596.000 775.010 600.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 596.000 74.890 600.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 596.000 125.030 600.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 596.000 175.170 600.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 596.000 224.850 600.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 596.000 274.990 600.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 596.000 325.130 600.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 596.000 375.270 600.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 596.000 424.950 600.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.810 596.000 475.090 600.000 ;
    END
  END io_oeb[9]
  PIN red[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.920 4.000 300.520 ;
    END
  END red[0]
  PIN red[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 385.600 4.000 386.200 ;
    END
  END red[1]
  PIN red[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.010 596.000 875.290 600.000 ;
    END
  END red[2]
  PIN red[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.960 4.000 557.560 ;
    END
  END red[3]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.560 4.000 129.160 ;
    END
  END reset
  PIN scl
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 74.840 900.000 75.440 ;
    END
  END scl
  PIN sda
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END sda
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 587.760 ;
    END
  END vssd1
  PIN vsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 224.440 900.000 225.040 ;
    END
  END vsync
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 894.240 587.605 ;
      LAYER met1 ;
        RECT 5.520 10.640 894.240 587.760 ;
      LAYER met2 ;
        RECT 7.450 595.720 24.650 596.770 ;
        RECT 25.490 595.720 74.330 596.770 ;
        RECT 75.170 595.720 124.470 596.770 ;
        RECT 125.310 595.720 174.610 596.770 ;
        RECT 175.450 595.720 224.290 596.770 ;
        RECT 225.130 595.720 274.430 596.770 ;
        RECT 275.270 595.720 324.570 596.770 ;
        RECT 325.410 595.720 374.710 596.770 ;
        RECT 375.550 595.720 424.390 596.770 ;
        RECT 425.230 595.720 474.530 596.770 ;
        RECT 475.370 595.720 524.670 596.770 ;
        RECT 525.510 595.720 574.350 596.770 ;
        RECT 575.190 595.720 624.490 596.770 ;
        RECT 625.330 595.720 674.630 596.770 ;
        RECT 675.470 595.720 724.770 596.770 ;
        RECT 725.610 595.720 774.450 596.770 ;
        RECT 775.290 595.720 824.590 596.770 ;
        RECT 825.430 595.720 874.730 596.770 ;
        RECT 875.570 595.720 890.470 596.770 ;
        RECT 7.450 4.280 890.470 595.720 ;
        RECT 7.450 4.000 74.790 4.280 ;
        RECT 75.630 4.000 224.750 4.280 ;
        RECT 225.590 4.000 374.710 4.280 ;
        RECT 375.550 4.000 524.670 4.280 ;
        RECT 525.510 4.000 674.630 4.280 ;
        RECT 675.470 4.000 824.590 4.280 ;
        RECT 825.430 4.000 890.470 4.280 ;
      LAYER met3 ;
        RECT 4.000 557.960 896.000 587.685 ;
        RECT 4.400 556.560 896.000 557.960 ;
        RECT 4.000 525.320 896.000 556.560 ;
        RECT 4.000 523.920 895.600 525.320 ;
        RECT 4.000 472.280 896.000 523.920 ;
        RECT 4.400 470.880 896.000 472.280 ;
        RECT 4.000 386.600 896.000 470.880 ;
        RECT 4.400 385.200 896.000 386.600 ;
        RECT 4.000 375.720 896.000 385.200 ;
        RECT 4.000 374.320 895.600 375.720 ;
        RECT 4.000 300.920 896.000 374.320 ;
        RECT 4.400 299.520 896.000 300.920 ;
        RECT 4.000 225.440 896.000 299.520 ;
        RECT 4.000 224.040 895.600 225.440 ;
        RECT 4.000 215.240 896.000 224.040 ;
        RECT 4.400 213.840 896.000 215.240 ;
        RECT 4.000 129.560 896.000 213.840 ;
        RECT 4.400 128.160 896.000 129.560 ;
        RECT 4.000 75.840 896.000 128.160 ;
        RECT 4.000 74.440 895.600 75.840 ;
        RECT 4.000 43.880 896.000 74.440 ;
        RECT 4.400 42.480 896.000 43.880 ;
        RECT 4.000 10.715 896.000 42.480 ;
      LAYER met4 ;
        RECT 281.815 11.735 327.840 371.105 ;
        RECT 330.240 11.735 404.640 371.105 ;
        RECT 407.040 11.735 481.440 371.105 ;
        RECT 483.840 11.735 494.665 371.105 ;
  END
END pong
END LIBRARY

