VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pong
  CLASS BLOCK ;
  FOREIGN pong ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN blue[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 596.000 750.170 600.000 ;
    END
  END blue[0]
  PIN blue[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 349.560 900.000 350.160 ;
    END
  END blue[1]
  PIN blue[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.210 0.000 562.490 4.000 ;
    END
  END blue[2]
  PIN blue[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 524.320 4.000 524.920 ;
    END
  END blue[3]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END clk
  PIN game_reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 49.680 900.000 50.280 ;
    END
  END game_reset
  PIN green[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.670 596.000 792.950 600.000 ;
    END
  END green[0]
  PIN green[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 449.520 900.000 450.120 ;
    END
  END green[1]
  PIN green[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.720 4.000 375.320 ;
    END
  END green[2]
  PIN green[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.230 596.000 878.510 600.000 ;
    END
  END green[3]
  PIN hsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END hsync
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 596.000 21.530 600.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 596.000 449.790 600.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 596.000 493.030 600.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 596.000 535.810 600.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 596.000 578.590 600.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.090 596.000 621.370 600.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 596.000 664.150 600.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 596.000 64.310 600.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 596.000 107.090 600.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 596.000 149.870 600.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 596.000 192.650 600.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 596.000 235.430 600.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 596.000 278.670 600.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 596.000 321.450 600.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 596.000 364.230 600.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.730 596.000 407.010 600.000 ;
    END
  END io_oeb[9]
  PIN red[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 249.600 900.000 250.200 ;
    END
  END red[0]
  PIN red[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.450 596.000 835.730 600.000 ;
    END
  END red[1]
  PIN red[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 549.480 900.000 550.080 ;
    END
  END red[2]
  PIN red[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.150 0.000 787.430 4.000 ;
    END
  END red[3]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END reset
  PIN scl
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.110 596.000 707.390 600.000 ;
    END
  END scl
  PIN sda
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 149.640 900.000 150.240 ;
    END
  END sda
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 587.760 ;
    END
  END vssd1
  PIN vsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END vsync
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 894.240 587.605 ;
      LAYER met1 ;
        RECT 5.520 10.640 894.240 587.760 ;
      LAYER met2 ;
        RECT 7.450 595.720 20.970 596.770 ;
        RECT 21.810 595.720 63.750 596.770 ;
        RECT 64.590 595.720 106.530 596.770 ;
        RECT 107.370 595.720 149.310 596.770 ;
        RECT 150.150 595.720 192.090 596.770 ;
        RECT 192.930 595.720 234.870 596.770 ;
        RECT 235.710 595.720 278.110 596.770 ;
        RECT 278.950 595.720 320.890 596.770 ;
        RECT 321.730 595.720 363.670 596.770 ;
        RECT 364.510 595.720 406.450 596.770 ;
        RECT 407.290 595.720 449.230 596.770 ;
        RECT 450.070 595.720 492.470 596.770 ;
        RECT 493.310 595.720 535.250 596.770 ;
        RECT 536.090 595.720 578.030 596.770 ;
        RECT 578.870 595.720 620.810 596.770 ;
        RECT 621.650 595.720 663.590 596.770 ;
        RECT 664.430 595.720 706.830 596.770 ;
        RECT 707.670 595.720 749.610 596.770 ;
        RECT 750.450 595.720 792.390 596.770 ;
        RECT 793.230 595.720 835.170 596.770 ;
        RECT 836.010 595.720 877.950 596.770 ;
        RECT 878.790 595.720 890.470 596.770 ;
        RECT 7.450 4.280 890.470 595.720 ;
        RECT 7.450 4.000 112.050 4.280 ;
        RECT 112.890 4.000 336.990 4.280 ;
        RECT 337.830 4.000 561.930 4.280 ;
        RECT 562.770 4.000 786.870 4.280 ;
        RECT 787.710 4.000 890.470 4.280 ;
      LAYER met3 ;
        RECT 4.000 550.480 896.000 587.685 ;
        RECT 4.000 549.080 895.600 550.480 ;
        RECT 4.000 525.320 896.000 549.080 ;
        RECT 4.400 523.920 896.000 525.320 ;
        RECT 4.000 450.520 896.000 523.920 ;
        RECT 4.000 449.120 895.600 450.520 ;
        RECT 4.000 375.720 896.000 449.120 ;
        RECT 4.400 374.320 896.000 375.720 ;
        RECT 4.000 350.560 896.000 374.320 ;
        RECT 4.000 349.160 895.600 350.560 ;
        RECT 4.000 250.600 896.000 349.160 ;
        RECT 4.000 249.200 895.600 250.600 ;
        RECT 4.000 225.440 896.000 249.200 ;
        RECT 4.400 224.040 896.000 225.440 ;
        RECT 4.000 150.640 896.000 224.040 ;
        RECT 4.000 149.240 895.600 150.640 ;
        RECT 4.000 75.840 896.000 149.240 ;
        RECT 4.400 74.440 896.000 75.840 ;
        RECT 4.000 50.680 896.000 74.440 ;
        RECT 4.000 49.280 895.600 50.680 ;
        RECT 4.000 10.715 896.000 49.280 ;
      LAYER met4 ;
        RECT 429.935 57.975 481.440 426.185 ;
        RECT 483.840 57.975 558.240 426.185 ;
        RECT 560.640 57.975 635.040 426.185 ;
        RECT 637.440 57.975 684.185 426.185 ;
  END
END pong
END LIBRARY

