magic
tech sky130A
magscale 1 2
timestamp 1653086684
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 2128 178848 117552
<< metal2 >>
rect 4250 119200 4306 120000
rect 12806 119200 12862 120000
rect 21362 119200 21418 120000
rect 29918 119200 29974 120000
rect 38474 119200 38530 120000
rect 47030 119200 47086 120000
rect 55678 119200 55734 120000
rect 64234 119200 64290 120000
rect 72790 119200 72846 120000
rect 81346 119200 81402 120000
rect 89902 119200 89958 120000
rect 98550 119200 98606 120000
rect 107106 119200 107162 120000
rect 115662 119200 115718 120000
rect 124218 119200 124274 120000
rect 132774 119200 132830 120000
rect 141422 119200 141478 120000
rect 149978 119200 150034 120000
rect 158534 119200 158590 120000
rect 167090 119200 167146 120000
rect 175646 119200 175702 120000
rect 22466 0 22522 800
rect 67454 0 67510 800
rect 112442 0 112498 800
rect 157430 0 157486 800
<< obsm2 >>
rect 1490 119144 4194 119354
rect 4362 119144 12750 119354
rect 12918 119144 21306 119354
rect 21474 119144 29862 119354
rect 30030 119144 38418 119354
rect 38586 119144 46974 119354
rect 47142 119144 55622 119354
rect 55790 119144 64178 119354
rect 64346 119144 72734 119354
rect 72902 119144 81290 119354
rect 81458 119144 89846 119354
rect 90014 119144 98494 119354
rect 98662 119144 107050 119354
rect 107218 119144 115606 119354
rect 115774 119144 124162 119354
rect 124330 119144 132718 119354
rect 132886 119144 141366 119354
rect 141534 119144 149922 119354
rect 150090 119144 158478 119354
rect 158646 119144 167034 119354
rect 167202 119144 175590 119354
rect 175758 119144 178094 119354
rect 1490 856 178094 119144
rect 1490 800 22410 856
rect 22578 800 67398 856
rect 67566 800 112386 856
rect 112554 800 157374 856
rect 157542 800 178094 856
<< metal3 >>
rect 179200 109896 180000 110016
rect 0 104864 800 104984
rect 179200 89904 180000 90024
rect 0 74944 800 75064
rect 179200 69912 180000 70032
rect 179200 49920 180000 50040
rect 0 44888 800 45008
rect 179200 29928 180000 30048
rect 0 14968 800 15088
rect 179200 9936 180000 10056
<< obsm3 >>
rect 800 110096 179200 117537
rect 800 109816 179120 110096
rect 800 105064 179200 109816
rect 880 104784 179200 105064
rect 800 90104 179200 104784
rect 800 89824 179120 90104
rect 800 75144 179200 89824
rect 880 74864 179200 75144
rect 800 70112 179200 74864
rect 800 69832 179120 70112
rect 800 50120 179200 69832
rect 800 49840 179120 50120
rect 800 45088 179200 49840
rect 880 44808 179200 45088
rect 800 30128 179200 44808
rect 800 29848 179120 30128
rect 800 15168 179200 29848
rect 880 14888 179200 15168
rect 800 10136 179200 14888
rect 800 9856 179120 10136
rect 800 2143 179200 9856
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 85987 11595 96288 85237
rect 96768 11595 111648 85237
rect 112128 11595 127008 85237
rect 127488 11595 136837 85237
<< labels >>
rlabel metal2 s 149978 119200 150034 120000 6 blue[0]
port 1 nsew signal output
rlabel metal3 s 179200 69912 180000 70032 6 blue[1]
port 2 nsew signal output
rlabel metal2 s 112442 0 112498 800 6 blue[2]
port 3 nsew signal output
rlabel metal3 s 0 104864 800 104984 6 blue[3]
port 4 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 clk
port 5 nsew signal input
rlabel metal3 s 179200 9936 180000 10056 6 game_reset
port 6 nsew signal input
rlabel metal2 s 158534 119200 158590 120000 6 green[0]
port 7 nsew signal output
rlabel metal3 s 179200 89904 180000 90024 6 green[1]
port 8 nsew signal output
rlabel metal3 s 0 74944 800 75064 6 green[2]
port 9 nsew signal output
rlabel metal2 s 175646 119200 175702 120000 6 green[3]
port 10 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 hsync
port 11 nsew signal output
rlabel metal2 s 4250 119200 4306 120000 6 io_oeb[0]
port 12 nsew signal output
rlabel metal2 s 89902 119200 89958 120000 6 io_oeb[10]
port 13 nsew signal output
rlabel metal2 s 98550 119200 98606 120000 6 io_oeb[11]
port 14 nsew signal output
rlabel metal2 s 107106 119200 107162 120000 6 io_oeb[12]
port 15 nsew signal output
rlabel metal2 s 115662 119200 115718 120000 6 io_oeb[13]
port 16 nsew signal output
rlabel metal2 s 124218 119200 124274 120000 6 io_oeb[14]
port 17 nsew signal output
rlabel metal2 s 132774 119200 132830 120000 6 io_oeb[15]
port 18 nsew signal output
rlabel metal2 s 12806 119200 12862 120000 6 io_oeb[1]
port 19 nsew signal output
rlabel metal2 s 21362 119200 21418 120000 6 io_oeb[2]
port 20 nsew signal output
rlabel metal2 s 29918 119200 29974 120000 6 io_oeb[3]
port 21 nsew signal output
rlabel metal2 s 38474 119200 38530 120000 6 io_oeb[4]
port 22 nsew signal output
rlabel metal2 s 47030 119200 47086 120000 6 io_oeb[5]
port 23 nsew signal output
rlabel metal2 s 55678 119200 55734 120000 6 io_oeb[6]
port 24 nsew signal output
rlabel metal2 s 64234 119200 64290 120000 6 io_oeb[7]
port 25 nsew signal output
rlabel metal2 s 72790 119200 72846 120000 6 io_oeb[8]
port 26 nsew signal output
rlabel metal2 s 81346 119200 81402 120000 6 io_oeb[9]
port 27 nsew signal output
rlabel metal3 s 179200 49920 180000 50040 6 red[0]
port 28 nsew signal output
rlabel metal2 s 167090 119200 167146 120000 6 red[1]
port 29 nsew signal output
rlabel metal3 s 179200 109896 180000 110016 6 red[2]
port 30 nsew signal output
rlabel metal2 s 157430 0 157486 800 6 red[3]
port 31 nsew signal output
rlabel metal2 s 67454 0 67510 800 6 reset
port 32 nsew signal input
rlabel metal2 s 141422 119200 141478 120000 6 scl
port 33 nsew signal bidirectional
rlabel metal3 s 179200 29928 180000 30048 6 sda
port 34 nsew signal bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 35 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 35 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 35 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 35 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 35 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 35 nsew power input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 36 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 36 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 36 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 36 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 36 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 36 nsew ground input
rlabel metal3 s 0 44888 800 45008 6 vsync
port 37 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 12871632
string GDS_FILE /home/debi/Desktop/Efabless_MFnJK/MPW6/mfNjK/pong-chip/openlane/pong/runs/pong/results/finishing/pong.magic.gds
string GDS_START 810400
<< end >>

