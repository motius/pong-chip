magic
tech sky130A
magscale 1 2
timestamp 1653069342
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 2128 178848 117552
<< metal2 >>
rect 4986 119200 5042 120000
rect 14922 119200 14978 120000
rect 24950 119200 25006 120000
rect 34978 119200 35034 120000
rect 44914 119200 44970 120000
rect 54942 119200 54998 120000
rect 64970 119200 65026 120000
rect 74998 119200 75054 120000
rect 84934 119200 84990 120000
rect 94962 119200 95018 120000
rect 104990 119200 105046 120000
rect 114926 119200 114982 120000
rect 124954 119200 125010 120000
rect 134982 119200 135038 120000
rect 145010 119200 145066 120000
rect 154946 119200 155002 120000
rect 164974 119200 165030 120000
rect 175002 119200 175058 120000
rect 15014 0 15070 800
rect 45006 0 45062 800
rect 74998 0 75054 800
rect 104990 0 105046 800
rect 134982 0 135038 800
rect 164974 0 165030 800
<< obsm2 >>
rect 1490 119144 4930 119354
rect 5098 119144 14866 119354
rect 15034 119144 24894 119354
rect 25062 119144 34922 119354
rect 35090 119144 44858 119354
rect 45026 119144 54886 119354
rect 55054 119144 64914 119354
rect 65082 119144 74942 119354
rect 75110 119144 84878 119354
rect 85046 119144 94906 119354
rect 95074 119144 104934 119354
rect 105102 119144 114870 119354
rect 115038 119144 124898 119354
rect 125066 119144 134926 119354
rect 135094 119144 144954 119354
rect 145122 119144 154890 119354
rect 155058 119144 164918 119354
rect 165086 119144 174946 119354
rect 175114 119144 178094 119354
rect 1490 856 178094 119144
rect 1490 800 14958 856
rect 15126 800 44950 856
rect 45118 800 74942 856
rect 75110 800 104934 856
rect 105102 800 134926 856
rect 135094 800 164918 856
rect 165086 800 178094 856
<< metal3 >>
rect 0 111392 800 111512
rect 179200 104864 180000 104984
rect 0 94256 800 94376
rect 0 77120 800 77240
rect 179200 74944 180000 75064
rect 0 59984 800 60104
rect 179200 44888 180000 45008
rect 0 42848 800 42968
rect 0 25712 800 25832
rect 179200 14968 180000 15088
rect 0 8576 800 8696
<< obsm3 >>
rect 800 111592 179200 117537
rect 880 111312 179200 111592
rect 800 105064 179200 111312
rect 800 104784 179120 105064
rect 800 94456 179200 104784
rect 880 94176 179200 94456
rect 800 77320 179200 94176
rect 880 77040 179200 77320
rect 800 75144 179200 77040
rect 800 74864 179120 75144
rect 800 60184 179200 74864
rect 880 59904 179200 60184
rect 800 45088 179200 59904
rect 800 44808 179120 45088
rect 800 43048 179200 44808
rect 880 42768 179200 43048
rect 800 25912 179200 42768
rect 880 25632 179200 25912
rect 800 15168 179200 25632
rect 800 14888 179120 15168
rect 800 8776 179200 14888
rect 880 8496 179200 8776
rect 800 2143 179200 8496
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 56363 2347 65568 74221
rect 66048 2347 80928 74221
rect 81408 2347 96288 74221
rect 96768 2347 98933 74221
<< labels >>
rlabel metal3 s 0 42848 800 42968 6 blue[0]
port 1 nsew signal output
rlabel metal3 s 179200 74944 180000 75064 6 blue[1]
port 2 nsew signal output
rlabel metal2 s 134982 0 135038 800 6 blue[2]
port 3 nsew signal output
rlabel metal2 s 164974 0 165030 800 6 blue[3]
port 4 nsew signal output
rlabel metal2 s 164974 119200 165030 120000 6 clk
port 5 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 game_reset
port 6 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 green[0]
port 7 nsew signal output
rlabel metal2 s 104990 0 105046 800 6 green[1]
port 8 nsew signal output
rlabel metal3 s 0 94256 800 94376 6 green[2]
port 9 nsew signal output
rlabel metal3 s 179200 104864 180000 104984 6 green[3]
port 10 nsew signal output
rlabel metal3 s 0 8576 800 8696 6 hsync
port 11 nsew signal output
rlabel metal2 s 4986 119200 5042 120000 6 io_oeb[0]
port 12 nsew signal output
rlabel metal2 s 104990 119200 105046 120000 6 io_oeb[10]
port 13 nsew signal output
rlabel metal2 s 114926 119200 114982 120000 6 io_oeb[11]
port 14 nsew signal output
rlabel metal2 s 124954 119200 125010 120000 6 io_oeb[12]
port 15 nsew signal output
rlabel metal2 s 134982 119200 135038 120000 6 io_oeb[13]
port 16 nsew signal output
rlabel metal2 s 145010 119200 145066 120000 6 io_oeb[14]
port 17 nsew signal output
rlabel metal2 s 154946 119200 155002 120000 6 io_oeb[15]
port 18 nsew signal output
rlabel metal2 s 14922 119200 14978 120000 6 io_oeb[1]
port 19 nsew signal output
rlabel metal2 s 24950 119200 25006 120000 6 io_oeb[2]
port 20 nsew signal output
rlabel metal2 s 34978 119200 35034 120000 6 io_oeb[3]
port 21 nsew signal output
rlabel metal2 s 44914 119200 44970 120000 6 io_oeb[4]
port 22 nsew signal output
rlabel metal2 s 54942 119200 54998 120000 6 io_oeb[5]
port 23 nsew signal output
rlabel metal2 s 64970 119200 65026 120000 6 io_oeb[6]
port 24 nsew signal output
rlabel metal2 s 74998 119200 75054 120000 6 io_oeb[7]
port 25 nsew signal output
rlabel metal2 s 84934 119200 84990 120000 6 io_oeb[8]
port 26 nsew signal output
rlabel metal2 s 94962 119200 95018 120000 6 io_oeb[9]
port 27 nsew signal output
rlabel metal3 s 0 59984 800 60104 6 red[0]
port 28 nsew signal output
rlabel metal3 s 0 77120 800 77240 6 red[1]
port 29 nsew signal output
rlabel metal2 s 175002 119200 175058 120000 6 red[2]
port 30 nsew signal output
rlabel metal3 s 0 111392 800 111512 6 red[3]
port 31 nsew signal output
rlabel metal3 s 0 25712 800 25832 6 reset
port 32 nsew signal input
rlabel metal3 s 179200 14968 180000 15088 6 scl
port 33 nsew signal bidirectional
rlabel metal2 s 45006 0 45062 800 6 sda
port 34 nsew signal bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 35 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 35 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 35 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 35 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 35 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 35 nsew power input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 36 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 36 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 36 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 36 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 36 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 36 nsew ground input
rlabel metal3 s 179200 44888 180000 45008 6 vsync
port 37 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 12883506
string GDS_FILE /home/debi/Desktop/Efabless_MFnJK/MPW6/mfNjK/pong-chip/openlane/pong/runs/pong/results/finishing/pong.magic.gds
string GDS_START 850122
<< end >>

